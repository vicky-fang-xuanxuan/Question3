/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  assign uio_out = 0;
  assign uio_oe  = 0;

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, clk, rst_n, 1'b0};

endmodule

module bitwise_majority (
    input  wire [7:0] A,      // First 8-bit input
    input  wire [7:0] B,      // Second 8-bit input
    output wire [7:0] C       // 8-bit Output
);

  assign C = (A & B) | (A ^ B); // Bitwise majority function

endmodule

module tb_bitwise_majority;
    reg [7:0] A, B;
    wire [7:0] C;

    bitwise_majority uut (
        .A(A),
        .B(B),
        .C(C)
    );

    initial begin
        $dumpfile("tb.vcd");
        $dumpvars(0, tb_bitwise_majority);

        // Test Cases
        A = 8'b11001100; B = 8'b10101010; #10;
        A = 8'b00000001; B = 8'b00000000; #10;
        A = 8'b11111111; B = 8'b00000000; #10;
        A = 8'b01010101; B = 8'b10101010; #10;

        $finish;
    end
endmodule
